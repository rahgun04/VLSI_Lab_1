##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Thu Oct  2 16:24:06 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO lfsr4
  CLASS BLOCK ;
  SIZE 17.400000 BY 17.000000 ;
  FOREIGN lfsr4 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 16.880000 7.650000 17.400000 7.750000 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 8.450000 0.520000 8.550000 ;
    END
  END rst
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.450000 16.480000 8.550000 17.000000 ;
    END
  END data_out[3]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.850000 16.480000 8.950000 17.000000 ;
    END
  END data_out[2]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.650000 0.000000 8.750000 0.520000 ;
    END
  END data_out[1]
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8.650000 0.000000 8.750000 0.520000 ;
    END
  END data_out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 17.400000 17.000000 ;
    LAYER M2 ;
      RECT 9.050000 16.380000 17.400000 17.000000 ;
      RECT 8.650000 16.380000 8.750000 17.000000 ;
      RECT 0.000000 16.380000 8.350000 17.000000 ;
      RECT 0.000000 0.620000 17.400000 16.380000 ;
      RECT 8.850000 0.000000 17.400000 0.620000 ;
      RECT 0.000000 0.000000 8.550000 0.620000 ;
    LAYER M3 ;
      RECT 0.000000 8.650000 17.400000 17.000000 ;
      RECT 0.620000 8.350000 17.400000 8.650000 ;
      RECT 0.000000 7.850000 17.400000 8.350000 ;
      RECT 0.000000 7.550000 16.780000 7.850000 ;
      RECT 0.000000 0.000000 17.400000 7.550000 ;
    LAYER M4 ;
      RECT 0.000000 0.620000 17.400000 17.000000 ;
      RECT 8.850000 0.000000 17.400000 0.620000 ;
      RECT 0.000000 0.000000 8.550000 0.620000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 17.400000 17.000000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 17.400000 17.000000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 17.400000 17.000000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 17.400000 17.000000 ;
    LAYER M9 ;
      RECT 0.000000 0.000000 17.400000 17.000000 ;
    LAYER AP ;
      RECT 0.000000 0.000000 17.400000 17.000000 ;
  END
END lfsr4

END LIBRARY
