##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Wed Oct  8 13:45:44 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO lfsr4
  CLASS BLOCK ;
  SIZE 46.400000 BY 11.400000 ;
  FOREIGN lfsr4 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.250000 10.880000 21.350000 11.400000 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.050000 10.880000 6.150000 11.400000 ;
    END
  END rst
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.050000 10.880000 33.150000 11.400000 ;
    END
  END data_out[3]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.050000 10.880000 28.150000 11.400000 ;
    END
  END data_out[2]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.250000 10.880000 13.350000 11.400000 ;
    END
  END data_out[1]
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.850000 10.880000 17.950000 11.400000 ;
    END
  END data_out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 46.400000 11.400000 ;
    LAYER M2 ;
      RECT 33.250000 10.780000 46.400000 11.400000 ;
      RECT 28.250000 10.780000 32.950000 11.400000 ;
      RECT 21.450000 10.780000 27.950000 11.400000 ;
      RECT 18.050000 10.780000 21.150000 11.400000 ;
      RECT 13.450000 10.780000 17.750000 11.400000 ;
      RECT 6.250000 10.780000 13.150000 11.400000 ;
      RECT 0.000000 10.780000 5.950000 11.400000 ;
      RECT 0.000000 0.000000 46.400000 10.780000 ;
    LAYER M3 ;
      RECT 0.000000 0.000000 46.400000 11.400000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 46.400000 11.400000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 46.400000 11.400000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 46.400000 11.400000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 46.400000 11.400000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 46.400000 11.400000 ;
    LAYER M9 ;
      RECT 0.000000 0.000000 46.400000 11.400000 ;
    LAYER AP ;
      RECT 0.000000 0.000000 46.400000 11.400000 ;
  END
END lfsr4

END LIBRARY
